module top(
    input clk,
    input reset
);

x1_8core CPU(clk, reset);

endmodule